
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity tb_CRCtransmitter is
end entity;

architecture sim of tb_CRCtransmitter is

    -- DUT signals
    signal clk         : std_logic := '0';
    signal input_data  : std_logic_vector(7 downto 0) := (others => '0');
    signal data_valid  : std_logic := '0';
    signal crc_out     : std_logic_vector(31 downto 0);

    -- Clock period
    constant CLK_PERIOD : time := 100 ps;

    -- ============================
    -- Test vector (EDIT HERE)
    -- ============================
    type byte_array is array (natural range <>) of std_logic_vector(7 downto 0);

    constant test_data : byte_array := ( --testing "ini ibu budi in ascii format" Bisa diganti sama data lain
       "01101001" , "01101110", "01101001", "00100000", "01101001", "01100010", "01110101", "00100000", "01100010", "01110101", "01100100", "01101001"

    );

begin

    -- ============================
    -- DUT instantiation
    -- ============================
    DUT : entity work.CRCtransmitter
        port map (
            input_data => input_data,
            crc_out    => crc_out,
            data_valid => data_valid,
            clk        => clk
        );

    -- ============================
    -- Clock generator
    -- ============================
    clk_process : process
    begin
        while true loop
            clk <= '0';
            wait for CLK_PERIOD / 2;
            clk <= '1';
            wait for CLK_PERIOD / 2;
        end loop;
    end process;

    -- ============================
    -- Stimulus process
    -- ============================
    stim_process : process
    begin
        -- Initial idle
        input_data <= (others => '0');
        data_valid <= '0';
        wait for CLK_PERIOD;

        -- Send bytes one per clock
        for i in test_data'range loop
            wait until rising_edge(clk);
            input_data <= test_data(i);
            data_valid <= '1';
        end loop;

        -- After last byte
        wait until rising_edge(clk);
        data_valid <= '0';
        input_data <= test_data(test_data'high); -- hold last value

        -- Stop simulation
        wait for 5 * CLK_PERIOD;
        assert false report "Simulation finished" severity failure;
    end process;

end architecture;