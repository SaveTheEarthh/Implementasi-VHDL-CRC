
-- Library
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Define entity
entity CRCreceiver is
	port	(
				input_data		:in		std_logic_vector (7 downto 0);	-- data A
                reset : in std_logic;
                data_valid  :in     std_logic;
				clk	:		in		std_logic;-- sinyal Clockian
                is_corrupt		: out  std_logic;
                crc_out		: out  STD_LOGIC_VECTOR(31 downto 0) -- data B -- data B
			);
end CRCreceiver;

-- Define architecture
architecture rtl of CRCreceiver is
    signal data_good, is_ready, is_4, en_regis: STD_LOGIC;
    signal  out_LUT1, out_LUT2, out_LUT3, out_LUT4, output_LUT, SIPO_out, data_after_regis32bit, data_after_XOR, data_after_LUT_prev: STD_LOGIC_VECTOR(31 downto 0);
    signal byteCount: STD_LOGIC_VECTOR(2 downto 0);
    signal first_byte, second_byte, third_byte, fourth_byte: STD_LOGIC_VECTOR(7 downto 0);
    signal padded_counter : std_logic_vector(31 downto 0);
signal padded_input   : std_logic_vector(31 downto 0);


component register32bitPIPO 
	port	(
			    A		:		in		std_logic_vector (31 downto 0);	-- data A
				En		:		in		std_logic;								-- sinyal Enable
				Res	    :		in		std_logic;								-- sinyal Reset
				Clk	    :		in		std_logic;								-- sinyal Clock
				Data	:		out	std_logic_vector (31 downto 0)		-- luaran data
			);
end component;

component Register32BitSIPO 
	port	(
        clk         : in  STD_LOGIC;
        reset       : in  STD_LOGIC;
        
        -- Interface ke UART (Input)
        uart_data   : in  STD_LOGIC_VECTOR (7 downto 0); -- Data 8-bit masuk
        uart_valid  : in  STD_LOGIC;                     -- Sinyal valid dari UART
        
        -- Interface ke CRC Engine (Output)
        chunk_data  : out STD_LOGIC_VECTOR (31 downto 0) -- Data 32-bit keluar      	-- luaran data
			);
end component;

component comparator 
	port	(
            inp_A,inp_B   : in std_logic_vector(31 downto 0);
	        equal : out std_logic
    );
end component;

component bytecounter 
	port	(
				clk             : in  STD_LOGIC;
                data_valid      : in  STD_LOGIC; -- Sinyal dari SIPO (Chunk Ready) -- Sinyal deteksi akhir (misal tombol/timeout)
        -- OUTPUT (Ke Datapath)
                currentCount    : out STD_LOGIC_VECTOR(2 downto 0)
			);
end component;

component CRC_Controller
  Port ( 
        -- INPUT (Dari Luar / Datapath)
        clk             : in  STD_LOGIC;
        is_4      : in  STD_LOGIC; -- Sinyal dari SIPO (Chunk Ready) -- Sinyal deteksi akhir (misal tombol/timeout)
        is_ready      : in  STD_LOGIC;
        -- OUTPUT (Ke Datapath)
        en_regis        : out STD_LOGIC -- Clock Enable Register -- Clock Enable Register
    );
end component;

component LUT_1
    Port ( addr_in : in  STD_LOGIC_VECTOR (7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (31 downto 0));
end component;

component LUT_2
Port ( addr_in : in  STD_LOGIC_VECTOR (7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (31 downto 0));
end component;

component LUT_3
Port ( addr_in : in  STD_LOGIC_VECTOR (7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (31 downto 0));
end component;

component LUT_4
Port ( addr_in : in  STD_LOGIC_VECTOR (7 downto 0);
           data_out : out  STD_LOGIC_VECTOR (31 downto 0));
end component;

component LUT_Prev
 Port ( 
        prev_crc_in : in  STD_LOGIC_VECTOR (31 downto 0); -- From Register
        lut_prev_out : out  STD_LOGIC_VECTOR (31 downto 0) -- To Feedback Mux/XOR
    );
end component;

begin

SIPO_atas: Register32BitSIPO
 port map(
    clk => clk,
    reset => reset,
    uart_data => input_data,
    uart_valid => data_valid,
    chunk_data => SIPO_out
);


CTRL: CRC_Controller
 port map(
    clk => clk,
    is_4 => is_4,
    is_ready => is_ready,
    en_regis => en_regis
);

first_byte <= SIPO_out(31 downto 24);
second_byte <= SIPO_out(23 downto 16);
third_byte <= SIPO_out(15 downto 8);
fourth_byte <= SIPO_out(7 downto 0);


LUT_1_inst: LUT_1
 port map(
    addr_in => first_byte,
    data_out => out_LUT1
);

LUT_2_inst: LUT_2
 port map(
    addr_in => second_byte,
    data_out => out_LUT2
);

LUT_3_inst: LUT_3
 port map(
    addr_in => third_byte,
    data_out => out_LUT3
);

LUT_4_inst: LUT_4
 port map(
    addr_in => fourth_byte,
    data_out => out_LUT4
);

LUT_Prev_inst: LUT_Prev
 port map(
    prev_crc_in => data_after_regis32bit,
    lut_prev_out => data_after_LUT_prev
);

output_LUT <= out_LUT1 xor out_LUT2 xor out_LUT3 xor out_LUT4;

data_after_XOR <= output_LUT xor data_after_LUT_prev;

-- Correct padding: 28 zeros + 4 bit counter = 32 bits
padded_counter <= "00000000000000000000000000000" & byteCount; 

-- Correct padding for input data check (checking against 32-bit comparator)
padded_input   <= "000000000000000000000000" & input_data;

REGIS_PIPO_bawah: register32bitPIPO
 port map(
    A => data_after_XOR,
    En => en_regis,
    Res => reset,
    Clk => Clk,
    Data => data_after_regis32bit
);

counter: byteCounter
	port map(
        Clk	=> Clk,
		data_valid	=> data_valid,
		currentCount => byteCount
	);

comparator_4: comparator
    port map(
        inp_A => padded_counter, -- Clean signal
        inp_B => "00000000000000000000000000000100",    -- Hex is cleaner than "000..100"
        equal => is_4
    );
comparator_ready: comparator
    port map(
        inp_A => padded_counter, -- Clean signal
        inp_B => "00000000000000000000000000000011",    -- Hex is cleaner than "000..100"
        equal => is_ready
    );

    crc_out <= data_after_regis32bit;

comparator_zero: comparator
    port map(
        inp_A => data_after_regis32bit, -- Clean signal
        inp_B => "00000000000000000000000000000000",    -- Hex is cleaner than "000..100"
        equal => data_good
    );
    is_corrupt <= not (data_good);

    end rtl;
	