library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
-- FSM oke, udah di simul sesuai
entity CRC_Controller is
    Port ( 
        -- INPUT (Dari Luar / Datapath)
        clk             : in  STD_LOGIC;
        is_4      : in  STD_LOGIC; -- Sinyal dari SIPO (Chunk Ready) -- Sinyal deteksi akhir (misal tombol/timeout)
        is_ready  :in  STD_LOGIC;

        -- OUTPUT (Ke Datapath)
        en_regis        : out STD_LOGIC -- Clock Enable Register-- Clock Enable Register
    );
end CRC_Controller;

architecture Behavioral of CRC_Controller is

    -- Definisi State
    type state_type is (
        S_IDLE,         -- Reset & Menunggu Data Pertama
        s_process,
        s_buffer   -- Menunggu SIPO penuh (4 byte pertama)         -- Selesai, Output Valid
    );
    
    signal current_state, next_state : state_type;

begin
    -- =========================================================
    -- PROSES 1: SEQUENTIAL (Memori State)
    -- =========================================================
    process(clk)
    begin
        if rising_edge(clk) then
            current_state <= next_state;
            end if;
           end process;

    -- =========================================================
    -- PROSES 2: COMBINATIONAL (Logika Transisi & Output)
    -- =========================================================
    process(current_state, is_4, is_ready)
    begin
        next_state <= current_state; -- Default stay

        case current_state is
            
            -- STATE: IDLE
            when S_IDLE =>
                en_regis <= '0'; -- Bersihkan SIPO
                -- Pindah ke tunggu data pertama
                if is_ready = '1' then
                    next_state <= s_buffer;
                else
                    next_state <= S_IDLE;
                end if;
            when s_buffer =>
                en_regis <= '1';
                if is_4 = '1' then
                    next_state <= s_process;
                else
                    next_state <= s_buffer;
                end if;
            -- STATE: MENUNGGU 4 BYTE PERTAMA
            when s_process =>
                en_regis <= '0'; -- Bersihkan SIPO
                -- Diam di sini sampai SIPO penuh
                if is_4 = '0' then
                    next_state <= S_IDLE;
                else
                    next_state <= S_IDLE;
                end if;

            
            -- STATE: MENUNGGU 4 BYTE SELANJUTNYA
           
        end case;
    end process;

end Behavioral;